*project netlist
.subckt NAND4 A B C E OUT VDD GND

M1 OUT A VDD VDD PCH L=65n W=200n
M2 OUT B VDD VDD PCH L=65n W=200n
M3 OUT C VDD VDD PCH L=65n W=200n
M4 OUT E VDD VDD PCH L=65n W=200n


M5 M5O E GND GND NCH L=65n W=200n
M6 M6O C M5O GND NCH L=65n W=200n
M7 M7O B M60 GND NCH L=65n W=200n
M8 MOUT A M7O GND NCH L=65n W=200n

.ends

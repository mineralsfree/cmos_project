*project netlist
.subckt NAND3 A B C OUT VDD GND

M1 OUT A VDD VDD PCH L=65n W=200n
M2 OUT B VDD VDD PCH L=65n W=200n
M3 OUT C VDD VDD PCH L=65n W=200n


M4 M4O C GND GND NCH L=65n W=200n
M5 M5O B M4O GND NCH L=65n W=200n
M6 OUT A M50 GND NCH L=65n W=200n

.ends

